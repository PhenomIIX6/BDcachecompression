module reqtestbench();
	logic [643:0] d;
	logic [63:0] tag;
	logic con, rd;
	logic [3:0] wordaddr;
	logic cachemiss;
	logic [643:0] deq;
	logic [63:0] taqeq;
	logic code110;
	requestfilter dut(.d(d), .tag(tag), .con(con), .wordaddr(wordaddr), .cachemiss(cachemiss));
	initial
		begin
			d = 644'b11010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010101010110; con = 1; tag = 64'hAAAAAAAAAAAAAAA0; rd = 1; wordaddr = 4'b0000; #40;
		end
endmodule