module testbench();
	logic [1087:0] readbuffer;
	logic [63:0] tag;
	logic con, clk, reset, rd, cachehit;
	logic [63:0] q;
	logic [3:0] addr;
	logic [3:0] wordaddr;
	logic [643:0] cq;
	logic [1023:0] dq;
	logic [643:0] cqic;
	cachewithcompression dut(.readbuffer(readbuffer), .tag(tag), .con(con), .clk(clk), .reset(reset), .rd(rd), .cachehit(cachehit));
	always
		begin
			clk = 1; #10; clk = 0; #10;
		end
	initial
		begin
			reset = 1; #80
			readbuffer = 1088'hAAAAAAAAAAAAAAA0ABCD0123DADA0000ABCD0123DADA1300ABCD0123DADA1488ABCD0123DADA1300ABCD0123DADA2323ABCD0123DADA1000ABCD0123DADA6666ABCD0123DADAFFFFABCD0123DADAAAAAABCD0123DADA1300ABCD0123DADA1300ABCD0123DADA1300ABCD0123DADA1300ABCD0123DADA1300ABCD0123DADA1300ABCD0123DADA1300; tag = 64'hAAAAAAAAAAAAAAAA; reset = 0; rd = 0; con = 1; #40;
			readbuffer = 1088'hAAAAAAAAAAAAAAA0ABCD0123DADA0000ABCD0123DADA1300ABCD0123DADA1488ABCD0123DADA1300ABCD0123DADA2323ABCD0123DADA1000ABCD0123DADA6666ABCD0123DADAFFFFABCD0123DADAAAAAABCD0123DADA1300ABCD0123DADA1300ABCD0123DADA1300ABCD0123DADA1300ABCD0123DADA1300ABCD0123DADA1300ABCD0123DADA1300; tag = 64'hAAAAAAAAAAAAAAAA; reset = 0; rd = 1; con = 1; #40;
		end
endmodule